** Profile: "2_ShutdownCurrent-2_ShutdownCurrent"  [ D:\1_WebUp\kakuninn\BD00C0A\TestCircuit\bd00c0awfp-pspicefiles\2_shutdowncurrent\2_shutdowncurrent.sim ] 

** Creating circuit file "2_ShutdownCurrent.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../bdxxc0axfp.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:

*Analysis directives: 
.DC LIN V_VCC 0 26.5 0.01 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\2_ShutdownCurrent.net" 


.END
